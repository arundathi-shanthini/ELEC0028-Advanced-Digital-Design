/*
Simple testbench file for com_struct.sv
Author: Arundathi Shaji Shanthini
*/

